<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-29.2882,2.49699,156.978,-104.436</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>12.5,-5.5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>21,-5.5</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>31,-5.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>40.5,-5</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>55.5,-5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>63.5,-5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>78,-5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>88,-5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>22,9</position>
<gparam>LABEL_TEXT BINARY ADDER (C=A+B)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_TOGGLE</type>
<position>12.5,-10.5</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>21.5,-10</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>30,-10</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_TOGGLE</type>
<position>39.5,-9.5</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_TOGGLE</type>
<position>55,-10</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_TOGGLE</type>
<position>66,-9.5</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_TOGGLE</type>
<position>78,-9</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>88,-9.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_FULLADDER_1BIT</type>
<position>83,-22.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_B_0</ID>27 </input>
<output>
<ID>OUT_0</ID>29 </output>
<input>
<ID>carry_in</ID>30 </input>
<output>
<ID>carry_out</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>98</ID>
<type>GA_LED</type>
<position>68.5,-44</position>
<input>
<ID>N_in2</ID>54 </input>
<input>
<ID>N_in3</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>GA_LED</type>
<position>54.5,-43.5</position>
<input>
<ID>N_in2</ID>55 </input>
<input>
<ID>N_in3</ID>34 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>GA_LED</type>
<position>40,-43</position>
<input>
<ID>N_in2</ID>57 </input>
<input>
<ID>N_in3</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>GA_LED</type>
<position>28.5,-43</position>
<input>
<ID>N_in2</ID>58 </input>
<input>
<ID>N_in3</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>67.5,-49.5</position>
<gparam>LABEL_TEXT C0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>54,-48.5</position>
<gparam>LABEL_TEXT C1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>40.5,-49</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>AA_LABEL</type>
<position>28.5,-49</position>
<gparam>LABEL_TEXT C3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>FF_GND</type>
<position>91.5,-25.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_FULLADDER_1BIT</type>
<position>58.5,-22</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_B_0</ID>31 </input>
<output>
<ID>OUT_0</ID>34 </output>
<input>
<ID>carry_in</ID>33 </input>
<output>
<ID>carry_out</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_FULLADDER_1BIT</type>
<position>36.5,-21.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_B_0</ID>37 </input>
<output>
<ID>OUT_0</ID>39 </output>
<input>
<ID>carry_in</ID>38 </input>
<output>
<ID>carry_out</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_FULLADDER_1BIT</type>
<position>17,-21</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_B_0</ID>41 </input>
<output>
<ID>OUT_0</ID>43 </output>
<input>
<ID>carry_in</ID>42 </input>
<output>
<ID>carry_out</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>121</ID>
<type>GA_LED</type>
<position>-3.5,-27</position>
<input>
<ID>N_in3</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>AA_TOGGLE</type>
<position>98.5,-17</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>103.5,-17</position>
<gparam>LABEL_TEXT SUB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>94.5,-64.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>55 </input>
<input>
<ID>IN_2</ID>57 </input>
<input>
<ID>IN_3</ID>58 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-19.5,82,-15.5</points>
<connection>
<GID>96</GID>
<name>IN_B_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>78,-15.5,78,-11</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>78,-15.5,82,-15.5</points>
<intersection>78 1</intersection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-19.5,84,-15.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>88,-15.5,88,-11.5</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>84,-15.5,88,-15.5</points>
<intersection>84 0</intersection>
<intersection>88 1</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-43,68.5,-34</points>
<connection>
<GID>98</GID>
<name>N_in3</name></connection>
<intersection>-34 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>83,-34,83,-25.5</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>68.5,-34,83,-34</points>
<intersection>68.5 0</intersection>
<intersection>83 1</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-24.5,91.5,-22.5</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-22.5,91.5,-22.5</points>
<connection>
<GID>96</GID>
<name>carry_in</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-19,57.5,-15.5</points>
<connection>
<GID>115</GID>
<name>IN_B_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>55,-15.5,55,-12</points>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>55,-15.5,57.5,-15.5</points>
<intersection>55 1</intersection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-19,59.5,-15.5</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>66,-15.5,66,-11.5</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59.5,-15.5,66,-15.5</points>
<intersection>59.5 0</intersection>
<intersection>66 1</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-22.5,70.5,-22</points>
<intersection>-22.5 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-22,70.5,-22</points>
<connection>
<GID>115</GID>
<name>carry_in</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-22.5,79,-22.5</points>
<connection>
<GID>96</GID>
<name>carry_out</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-42.5,54.5,-33.5</points>
<connection>
<GID>100</GID>
<name>N_in3</name></connection>
<intersection>-33.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>58.5,-33.5,58.5,-25</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<intersection>-33.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-33.5,58.5,-33.5</points>
<intersection>54.5 0</intersection>
<intersection>58.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,-26,-3.5,-21</points>
<connection>
<GID>121</GID>
<name>N_in3</name></connection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3.5,-21,13,-21</points>
<connection>
<GID>119</GID>
<name>carry_out</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-18.5,37.5,-15</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>39.5,-15,39.5,-11.5</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-15,39.5,-15</points>
<intersection>37.5 0</intersection>
<intersection>39.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-18.5,35.5,-15</points>
<connection>
<GID>117</GID>
<name>IN_B_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>30,-15,30,-12</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30,-15,35.5,-15</points>
<intersection>30 1</intersection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-22,47.5,-21.5</points>
<intersection>-22 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-21.5,47.5,-21.5</points>
<connection>
<GID>117</GID>
<name>carry_in</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47.5,-22,54.5,-22</points>
<connection>
<GID>115</GID>
<name>carry_out</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-42,40,-33</points>
<connection>
<GID>102</GID>
<name>N_in3</name></connection>
<intersection>-33 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>36.5,-33,36.5,-24.5</points>
<connection>
<GID>117</GID>
<name>OUT_0</name></connection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-33,40,-33</points>
<intersection>36.5 1</intersection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-18,18,-15</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>21.5,-15,21.5,-12</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>18,-15,21.5,-15</points>
<intersection>18 0</intersection>
<intersection>21.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-18,16,-15</points>
<connection>
<GID>119</GID>
<name>IN_B_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>12.5,-15,12.5,-12.5</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-15,16,-15</points>
<intersection>12.5 1</intersection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-21.5,26.5,-21</points>
<intersection>-21.5 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-21,26.5,-21</points>
<connection>
<GID>119</GID>
<name>carry_in</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-21.5,32.5,-21.5</points>
<connection>
<GID>117</GID>
<name>carry_out</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-42,28.5,-33</points>
<connection>
<GID>104</GID>
<name>N_in3</name></connection>
<intersection>-33 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>17,-33,17,-24</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>17,-33,28.5,-33</points>
<intersection>17 1</intersection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-67.5,68.5,-45</points>
<connection>
<GID>98</GID>
<name>N_in2</name></connection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-67.5,89.5,-67.5</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-66.5,54.5,-44.5</points>
<connection>
<GID>100</GID>
<name>N_in2</name></connection>
<intersection>-66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-66.5,89.5,-66.5</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-65.5,40,-44</points>
<connection>
<GID>102</GID>
<name>N_in2</name></connection>
<intersection>-65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-65.5,89.5,-65.5</points>
<connection>
<GID>144</GID>
<name>IN_2</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-64.5,28.5,-44</points>
<connection>
<GID>104</GID>
<name>N_in2</name></connection>
<intersection>-64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-64.5,89.5,-64.5</points>
<connection>
<GID>144</GID>
<name>IN_3</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-23.2667,13.3667,163,-93.5667</PageViewport>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>17,-5</position>
<gparam>LABEL_TEXT HALF ADDER</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>15.5,-12.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>15.5,-21.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_AND2</type>
<position>37.5,-14.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AI_XOR2</type>
<position>38,-24</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>20.5,-13</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>20.5,-21.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>31</ID>
<type>HE_JUNC_4</type>
<position>25,-13</position>
<input>
<ID>N_in0</ID>1 </input>
<input>
<ID>N_in1</ID>6 </input>
<input>
<ID>N_in3</ID>3 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>HE_JUNC_4</type>
<position>24.5,-21.5</position>
<input>
<ID>N_in0</ID>2 </input>
<input>
<ID>N_in1</ID>5 </input>
<input>
<ID>N_in3</ID>4 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>45,-14.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>GA_LED</type>
<position>45,-24</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>51,-23.5</position>
<gparam>LABEL_TEXT SUM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>52.5,-14</position>
<gparam>LABEL_TEXT CARRY</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>18,-31</position>
<gparam>LABEL_TEXT FULL ADDER</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>15.5,-43</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>15,-54</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>15.5,-67</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>55.5,-31.5</position>
<gparam>LABEL_TEXT SUM = A XOR B XOR C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>54.5,-35.5</position>
<gparam>LABEL_TEXT CARRY= AB+AC+BC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>21.5,-43</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_TOGGLE</type>
<position>21,-55</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_TOGGLE</type>
<position>20,-67</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>HE_JUNC_4</type>
<position>26.5,-43.5</position>
<input>
<ID>N_in0</ID>9 </input>
<input>
<ID>N_in1</ID>16 </input>
<input>
<ID>N_in2</ID>18 </input>
<input>
<ID>N_in3</ID>12 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>HE_JUNC_4</type>
<position>26.5,-55</position>
<input>
<ID>N_in0</ID>10 </input>
<input>
<ID>N_in1</ID>17 </input>
<input>
<ID>N_in2</ID>20 </input>
<input>
<ID>N_in3</ID>13 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>HE_JUNC_4</type>
<position>26,-67</position>
<input>
<ID>N_in0</ID>11 </input>
<input>
<ID>N_in1</ID>19 </input>
<input>
<ID>N_in2</ID>21 </input>
<input>
<ID>N_in3</ID>14 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AI_XOR3</type>
<position>47,-69.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<input>
<ID>IN_2</ID>14 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>64</ID>
<type>GA_LED</type>
<position>55,-69.5</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>61,-69</position>
<gparam>LABEL_TEXT SUM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_AND2</type>
<position>47.5,-43.5</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_AND2</type>
<position>47.5,-49.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_AND2</type>
<position>47.5,-56</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>AE_OR3</type>
<position>60,-48.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>23 </input>
<input>
<ID>IN_2</ID>24 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>75</ID>
<type>GA_LED</type>
<position>68,-48.5</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>78.5,-48.5</position>
<gparam>LABEL_TEXT CARRY</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-13,24,-13</points>
<connection>
<GID>31</GID>
<name>N_in0</name></connection>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-21.5,23.5,-21.5</points>
<connection>
<GID>33</GID>
<name>N_in0</name></connection>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-12,25,-11</points>
<connection>
<GID>31</GID>
<name>N_in3</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-11,34.5,-11</points>
<intersection>25 0</intersection>
<intersection>34.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>34.5,-13.5,34.5,-11</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-11 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-20.5,24.5,-15.5</points>
<connection>
<GID>33</GID>
<name>N_in3</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-15.5,34.5,-15.5</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-23,30,-21.5</points>
<intersection>-23 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-23,35,-23</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-21.5,30,-21.5</points>
<connection>
<GID>33</GID>
<name>N_in1</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-25,30.5,-13</points>
<intersection>-25 1</intersection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-25,35,-25</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-13,30.5,-13</points>
<connection>
<GID>31</GID>
<name>N_in1</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-14.5,44,-14.5</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<connection>
<GID>35</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-24,44,-24</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<connection>
<GID>37</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23.5,-43,25.5,-43</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>25.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25.5,-43.5,25.5,-43</points>
<connection>
<GID>56</GID>
<name>N_in0</name></connection>
<intersection>-43 1</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-55,25.5,-55</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>25.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>25.5,-55,25.5,-55</points>
<connection>
<GID>58</GID>
<name>N_in0</name></connection>
<intersection>-55 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-67,25,-67</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<connection>
<GID>60</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-67.5,32.5,-42.5</points>
<intersection>-67.5 1</intersection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-67.5,44,-67.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-42.5,32.5,-42.5</points>
<connection>
<GID>56</GID>
<name>N_in3</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-69.5,29.5,-54</points>
<intersection>-69.5 1</intersection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-69.5,44,-69.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-54,29.5,-54</points>
<connection>
<GID>58</GID>
<name>N_in3</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-71.5,28,-66</points>
<intersection>-71.5 1</intersection>
<intersection>-66 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-71.5,44,-71.5</points>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-66,28,-66</points>
<connection>
<GID>60</GID>
<name>N_in3</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-69.5,54,-69.5</points>
<connection>
<GID>64</GID>
<name>N_in0</name></connection>
<connection>
<GID>62</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-43.5,36,-42.5</points>
<intersection>-43.5 2</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-42.5,44.5,-42.5</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-43.5,36,-43.5</points>
<connection>
<GID>56</GID>
<name>N_in1</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-55,36,-44.5</points>
<intersection>-55 2</intersection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-44.5,44.5,-44.5</points>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-55,36,-55</points>
<connection>
<GID>58</GID>
<name>N_in1</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-48.5,26.5,-44.5</points>
<connection>
<GID>56</GID>
<name>N_in2</name></connection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-48.5,44.5,-48.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-67,35.5,-50.5</points>
<intersection>-67 2</intersection>
<intersection>-50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-50.5,44.5,-50.5</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-67,35.5,-67</points>
<connection>
<GID>60</GID>
<name>N_in1</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-56,26.5,-55</points>
<connection>
<GID>58</GID>
<name>N_in2</name></connection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-55,44.5,-55</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-68,26,-57</points>
<connection>
<GID>60</GID>
<name>N_in2</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-57,44.5,-57</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-46.5,53.5,-43.5</points>
<intersection>-46.5 1</intersection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-46.5,57,-46.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-43.5,53.5,-43.5</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-49.5,53.5,-48.5</points>
<intersection>-49.5 2</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-48.5,57,-48.5</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-49.5,53.5,-49.5</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-56,53.5,-50.5</points>
<intersection>-56 2</intersection>
<intersection>-50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-50.5,57,-50.5</points>
<connection>
<GID>73</GID>
<name>IN_2</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-56,53.5,-56</points>
<connection>
<GID>71</GID>
<name>OUT</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,-48.5,67,-48.5</points>
<connection>
<GID>75</GID>
<name>N_in0</name></connection>
<connection>
<GID>73</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,0,139.7,-80.2</PageViewport>
<gate>
<ID>129</ID>
<type>AA_LABEL</type>
<position>22.5,-4</position>
<gparam>LABEL_TEXT ONES Complement</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>131</ID>
<type>AA_LABEL</type>
<position>18.5,-12.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_LABEL</type>
<position>45,-25</position>
<gparam>LABEL_TEXT SUB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>134</ID>
<type>AA_TOGGLE</type>
<position>18,-18</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>136</ID>
<type>AA_TOGGLE</type>
<position>40,-25</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>138</ID>
<type>AI_XOR2</type>
<position>22.5,-34</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>140</ID>
<type>GA_LED</type>
<position>22.5,-48.5</position>
<input>
<ID>N_in3</ID>52 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>AA_LABEL</type>
<position>30.5,-49</position>
<gparam>LABEL_TEXT ~B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-31,23.5,-25</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-25,38,-25</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-31,21.5,-25.5</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>18,-25.5,18,-20</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>18,-25.5,21.5,-25.5</points>
<intersection>18 1</intersection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-47.5,22.5,-37</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<connection>
<GID>140</GID>
<name>N_in3</name></connection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,0,139.7,-80.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.7,-80.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.7,-80.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.7,-80.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.7,-80.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.7,-80.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.7,-80.2</PageViewport></page 9></circuit>